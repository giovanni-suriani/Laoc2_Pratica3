module unidade_despacho(
    input Clock, 
    input Reset, 
    output Instrucao_i, 
    output Instrucao_l);
endmodule