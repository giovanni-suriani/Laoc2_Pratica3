module estacao_reserva_l(
    input Clock,
    input [15:0] Instrucao,
    input Reset
);
endmodule