module CDB_arbiter (
  input Clock,
  input Reset,
  output [15:0] CDB
);

endmodule