module CDB(
    input Reset, 
    input Estacao_i_out,
    input Estacao_l_out
);

endmodule