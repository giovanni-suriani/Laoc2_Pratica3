module tomasulo(input Clock,
                    input Reset);
                    
endmodule
