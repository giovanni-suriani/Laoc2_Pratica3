module CDB_arbiter (
  input Clock,
  input Reset,
  output reg [2:0]  Qi_CDB,
  output reg [15:0] Qi_CDB_Data
);

endmodule